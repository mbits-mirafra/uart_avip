
`ifndef UARTRxSEQUENCEPKG_INCLUDED_
`define UARTRxSEQUENCEPKG_INCLUDED_

package UartRxSequencePkg;
  import uvm_pkg :: *;
  `include "uvm_macros.svh"
  import UartGlobalPkg :: *;
  import UartRxPkg ::*;

  `include"UartRxBaseSequence.sv"
 
endpackage
`endif
